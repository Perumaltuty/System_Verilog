`timescale 1ns / 1ps
module repeat_for;
initial begin
  for (int i = 1;i<=4;i++)begin  
    $display ("Smart");   
    $display ("IOPS");
    end 
end 
endmodule 
